`include "baseclass.sv"
`include "transaction.sv"
`include "interface.sv"
`define Ntimes 50000
