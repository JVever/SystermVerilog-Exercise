interface alu_if;
	logic [3:0] a, b;
	logic [2:0] select;
	logic [4:0] result;
endinterface
